module control_unit(

input clk,
input N_flag,
input lsb,
input [8:0] addr, //first 9 bit of micro instruction
input [8:0] IR, //opcode in IR
output reg [35:0] MIR

);

reg [35:0] ROM[0:75]; // 76 micro instructions and 36bit length control signals

reg [3:0] mux_sel;
// parameter define
parameter FETCH4 = 9'd3;
parameter JUMPLSB = 9'd63;
parameter JUMPNLSB = 9'd67;
parameter JUMPNEG = 9'd71;

parameter STORER3 = 9'd24;

parameter LDARC3 = 9'd13;
parameter LOAD3 = 9'd20;
parameter STACR3 = 9'd27;
parameter ADD3 = 9'd44;
parameter MULR3 = 9'd61;
parameter SUB3 = 9'd48;


parameter
Rcol = 9'b000000001,
Rrow = 9'b000000010,
Ri   = 9'b000000011, 
Rj   = 9'b000000100, 
Rtotal = 9'b000000101, 
Raddress = 9'b000000110, 
Rbnd  = 9'b000000111, 
RcolTemp = 9'b000001000;

parameter
rcol_sel = 4'b0011,
rrow_sel = 4'b0100,
ri_sel   = 4'b0101,
rj_sel   = 4'b0110,
rtotal_sel   = 4'b0111,
raddress_sel = 4'b1000,
rbnd_sel     = 4'b1001,
rcoltemp_sel = 4'b1010;

initial 
	begin
		MIR = 36'b0;

	end


always @(negedge clk)
begin
    mux_sel =   (IR == Rcol)? rcol_sel :
                (IR == Rrow)? rrow_sel :
                (IR == Ri)? ri_sel :
                (IR == Rj)? rj_sel :
                (IR == Rtotal)? rtotal_sel :
                (IR == Raddress)? raddress_sel :
                (IR == Rbnd)? rbnd_sel :
                (IR == RcolTemp)? rcoltemp_sel:  4'b0;
                
        case(addr)
            FETCH4 : MIR = {IR,ROM[FETCH4][26:0]};

            JUMPLSB  : if (lsb == 1'b0) MIR = {9'd64,ROM[JUMPLSB][26:0]};
                        else MIR = {9'd66,ROM[JUMPLSB][26:0]};
            
            JUMPNLSB  : if (lsb == 1'b1) MIR = {9'd68,ROM[JUMPNLSB][26:0]};
                        else MIR = {9'd70,ROM[JUMPNLSB][26:0]};

            JUMPNEG  : if (N_flag == 1'b1) MIR = {9'd72,ROM[JUMPNEG][26:0]};
                       else MIR = {9'd74,ROM[JUMPNEG][26:0]};         

            STORER3  : MIR = {ROM[STORER3][35:18],IR[3:0],ROM[STORER3][13:0]};

            LDARC3 :  MIR = {ROM[LDARC3][35:7],mux_sel,ROM[LDARC3][2:0]};
            LOAD3  :  MIR = {ROM[LOAD3][35:7],mux_sel,ROM[LOAD3][2:0]};
            STACR3 :  MIR = {ROM[STACR3][35:7],mux_sel,ROM[STACR3][2:0]};
            ADD3   :  MIR = {ROM[ADD3][35:7],mux_sel,ROM[ADD3][2:0]};
            MULR3  :  MIR = {ROM[MULR3][35:7],mux_sel,ROM[MULR3][2:0]};
            SUB3   :  MIR = {ROM[SUB3][35:7],mux_sel,ROM[SUB3][2:0]};

            default : MIR = ROM[addr];


        endcase
	end
// define the microinstruction in the control store
initial 
begin

ROM[0] =36'b000000001_010000000_0000_0_00_0000_0000_00_0;
ROM[1] =36'b000000010_000000001_0000_0_01_0000_0000_00_0;
ROM[2] =36'b000000011_010100000_0000_0_00_0000_0000_00_0;
ROM[3] =36'bXXXXXXXXX_000000000_0000_0_00_0000_0000_00_0;

ROM[4] =36'b000000101_000000001_0000_0_11_0000_0000_00_0;
ROM[5] =36'b000000110_001000001_0000_0_01_0000_0000_00_0;
ROM[6] =36'b000000111_000000000_0000_0_00_1101_0001_01_0;
ROM[7] =36'b000001000_000010000_0000_0_00_0000_0000_00_0;
ROM[8] =36'b000001001_000001000_0000_0_00_0000_0000_00_0;
ROM[9] =36'b000001010_000000000_0000_0_00_0001_0010_00_0;
ROM[10]=36'b000000000_000000010_0000_0_00_0000_0000_00_0;

ROM[11]=36'b000001100_000000001_0000_0_01_0000_0000_00_0;
ROM[12]=36'b000001101_000100000_0000_0_00_0000_0000_00_0;
ROM[13]=36'b000001110_000000000_0000_0_00_0001_XXXX_00_0;
ROM[14]=36'b000001111_000010000_0000_0_00_0000_0000_00_0;
ROM[15]=36'b000010000_000001000_0000_0_00_0000_0000_00_0;
ROM[16]=36'b000010001_000000000_0000_0_00_0001_0000_00_0;
ROM[17]=36'b000000000_000000010_0000_0_00_0000_0000_00_0;

ROM[18]=36'b000010011_000000001_0000_0_01_0000_0000_00_0;
ROM[19]=36'b000010100_000100000_0000_0_00_0000_0000_00_0;
ROM[20]=36'b000010101_000000000_0000_0_00_0001_XXXX_00_0;
ROM[21]=36'b000000000_000000010_0000_0_00_0000_0000_00_0;

ROM[22]=36'b000010111_000000001_0000_0_01_0010_0000_10_0;
ROM[23]=36'b000011000_000100000_0000_0_00_0000_0000_00_0;
ROM[24]=36'b000000000_000000000_0000_0_00_0000_0000_00_0;

ROM[25]=36'b000011010_000000001_0000_0_01_0010_0000_10_0;
ROM[26]=36'b000011011_000100100_0000_0_00_0000_0000_00_0;
ROM[27]=36'b000011100_000000000_0000_0_00_0001_XXXX_00_0;
ROM[28]=36'b000011101_000010000_0000_0_00_0000_0000_00_0;
ROM[29]=36'b000000000_000000000_0000_1_00_0000_0000_00_0;

ROM[30]=36'b000011111_000000000_0000_0_00_0011_0000_10_0;
ROM[31]=36'b000000000_000000010_0000_0_00_0000_0000_00_0;

ROM[32]=36'b000100001_000000000_0000_0_00_0100_0000_10_0;
ROM[33]=36'b000000000_000000010_0000_0_00_0000_0000_00_0;

ROM[34]=36'b000100011_000000000_0000_0_00_0101_0000_10_0;
ROM[35]=36'b000000000_000000010_0000_0_00_0000_0000_00_0;

ROM[36]=36'b000100101_000000000_0000_0_00_0110_0000_10_0;
ROM[37]=36'b000000000_000000010_0000_0_00_0000_0000_00_0;

ROM[38]=36'b000100111_000000000_0000_0_00_0111_0000_10_0;
ROM[39]=36'b000000000_000000010_0000_0_00_0000_0000_00_0;

ROM[40]=36'b000101001_000000000_0000_0_00_1000_0000_10_0;
ROM[41]=36'b000000000_000000010_0000_0_00_0000_0000_00_0;

ROM[42]=36'b000101011_000000001_0000_0_01_0000_0000_00_0;
ROM[43]=36'b000101100_000100000_0000_0_00_0000_0000_00_0;
ROM[44]=36'b000101101_000000000_0000_0_00_1001_XXXX_10_0;
ROM[45]=36'b000000000_000000010_0000_0_00_0000_0000_00_0;

ROM[46]=36'b000101111_000000001_0000_0_01_0000_0000_00_0;
ROM[47]=36'b000110000_000100000_0000_0_00_0000_0000_00_0;
ROM[48]=36'b000110001_000000000_0000_0_00_1010_XXXX_10_0;
ROM[49]=36'b000000000_000000010_0000_0_00_0000_0000_00_0;

ROM[50]=36'b000110011_000000001_0000_0_01_0000_0000_00_0;
ROM[51]=36'b000110100_000000000_0000_0_00_1011_0001_10_0;
ROM[52]=36'b000000000_000000010_0000_0_00_0000_0000_00_0;

ROM[53]=36'b000110110_000000001_0000_0_01_0000_0000_00_0;
ROM[54]=36'b000110111_000000000_0000_0_00_1100_0001_10_0;
ROM[55]=36'b000000000_000000010_0000_0_00_0000_0000_00_0;

ROM[56]=36'b000111001_000000001_0000_0_01_0000_0000_00_0;
ROM[57]=36'b000111010_000000000_0000_0_00_0001_0001_00_0;
ROM[58]=36'b000000000_000000010_0000_0_00_0000_0000_00_0;

ROM[59]=36'b000111100_000000001_0000_0_01_0000_0000_00_0;
ROM[60]=36'b000111101_000100000_0000_0_00_0000_0000_00_0;
ROM[61]=36'b000111110_000000000_0000_0_00_1011_XXXX_10_0;
ROM[62]=36'b000000000_000000010_0000_0_00_0000_0000_00_0;

ROM[63]=36'bXXXXXXXXX_000000000_0000_0_00_0000_0000_00_0;
ROM[64]=36'b001000001_000000001_0000_0_00_0000_0000_00_0;
ROM[65]=36'b000000000_100000000_0000_0_00_0000_0000_00_0;
ROM[66]=36'b000000000_000000000_0000_0_01_0000_0000_00_0;

ROM[67]=36'bXXXXXXXXX_000000000_0000_0_00_0000_0000_00_0;
ROM[68]=36'b001000101_000000001_0000_0_00_0000_0000_00_0;
ROM[69]=36'b000000000_100000000_0000_0_00_0000_0000_00_0;
ROM[70]=36'b000000000_000000000_0000_0_01_0000_0000_00_0;

ROM[71]=36'bXXXXXXXXX_000000000_0000_0_00_0000_0000_00_0;
ROM[72]=36'b001001001_000000001_0000_0_00_0000_0000_00_0;
ROM[73]=36'b000000000_100000000_0000_0_00_0000_0000_00_0;
ROM[74]=36'b000000000_000000000_0000_0_01_0000_0000_00_0;

ROM[75]=36'bXXXXXXXXX_000000000_0000_0_01_0000_0000_00_1;


end
endmodule
